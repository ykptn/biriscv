module tb_poly_horner_mul;

reg clk;
reg rst;

localparam PASS_PC = 32'h80000130;
localparam FAIL_PC = 32'h80000134;
localparam UART_BASE = 32'h9200_0000;
localparam UART_SHADOW_ADDR = 32'h80018000;

reg [7:0] mem[131072:0];
integer i;
integer f;

initial begin
    $display("Starting POLY HORNER MUL EDP benchmark");

    if (`TRACE) begin
        $dumpfile("waveform.vcd");
        $dumpvars(0, tb_poly_horner_mul);
    end

    clk = 0;
    rst = 1;
    repeat (5) @(posedge clk);
    rst = 0;

    for (i = 0; i < 131072; i = i + 1)
        mem[i] = 0;

    f = $fopenr("./build/tcm.bin");
    i = $fread(mem, f);
    $display("Loaded %0d bytes from tcm.bin", i);
    for (i = 0; i < 131072; i = i + 1)
        u_mem.write(i, mem[i]);

    $display("RAM[0] = 0x%016h", u_mem.u_ram.ram[0]);
    $display("RAM[1] = 0x%016h", u_mem.u_ram.ram[1]);
    $display("RAM[2] = 0x%016h", u_mem.u_ram.ram[2]);
end

reg [63:0] cycle_count;
reg pass_reported;
reg fail_reported;
reg pass_pending;
reg [3:0] pass_delay;

initial begin
    cycle_count   = 0;
    pass_reported = 1'b0;
    fail_reported = 1'b0;
    pass_pending  = 1'b0;
    pass_delay    = 4'd0;
end

always @(posedge clk) begin
    if (rst) begin
        cycle_count   <= 0;
        pass_reported <= 1'b0;
        fail_reported <= 1'b0;
        pass_pending  <= 1'b0;
        pass_delay    <= 4'd0;
    end else begin
        cycle_count <= cycle_count + 1;

        if (!pass_pending && mem_i_pc_w == PASS_PC)
        begin
            pass_pending <= 1'b1;
            pass_delay   <= 4'd8;
        end
        else if (pass_pending && pass_delay != 0)
            pass_delay <= pass_delay - 1'b1;

        if (pass_pending && pass_delay == 0 && !pass_reported)
        begin
            pass_reported <= 1'b1;
            $display("\n*** POLY HORNER MUL EDP PASS ***");
            $finish;
        end
        else if (!fail_reported && mem_i_pc_w == FAIL_PC)
        begin
            fail_reported <= 1'b1;
            $display("\n*** POLY HORNER MUL EDP FAIL ***");
            $finish;
        end
        else if (cycle_count > 200000 && !pass_reported && !fail_reported)
        begin
            fail_reported <= 1'b1;
            $display("\nTimeout after %0d cycles (last PC 0x%08h)", cycle_count, mem_i_pc_w);
            $finish;
        end
    end
end

wire uart_write_w = (mem_d_wr_w != 4'b0) && (mem_d_addr_w == UART_BASE);

always @(posedge clk) begin
    if (!rst && uart_write_w) begin
        $write("%c", mem_d_data_wr_w[7:0]);
    end
end

initial begin
    forever clk = #5 ~clk;
end

wire          mem_i_rd_w;
wire          mem_i_flush_w;
wire          mem_i_invalidate_w;
wire [ 31:0]  mem_i_pc_w;
wire [ 31:0]  mem_d_addr_w;
wire [ 31:0]  mem_d_data_wr_w;
wire          mem_d_rd_w;
wire [  3:0]  mem_d_wr_w;
wire          mem_d_cacheable_w;
wire [ 10:0]  mem_d_req_tag_w;
wire          mem_d_invalidate_w;
wire          mem_d_writeback_w;
wire          mem_d_flush_w;
wire          mem_i_accept_w;
wire          mem_i_valid_w;
wire          mem_i_error_w;
wire [ 63:0]  mem_i_inst_w;
wire [ 31:0]  mem_d_data_rd_w;
wire          mem_d_accept_w;
wire          mem_d_ack_w;
wire          mem_d_error_w;
wire [ 10:0]  mem_d_resp_tag_w;

wire [31:0] mem_d_addr_mem_w = uart_write_w ? UART_SHADOW_ADDR : mem_d_addr_w;

riscv_core u_dut
(
     .clk_i(clk)
    ,.rst_i(rst)
    ,.mem_d_data_rd_i(mem_d_data_rd_w)
    ,.mem_d_accept_i(mem_d_accept_w)
    ,.mem_d_ack_i(mem_d_ack_w)
    ,.mem_d_error_i(mem_d_error_w)
    ,.mem_d_resp_tag_i(mem_d_resp_tag_w)
    ,.mem_i_accept_i(mem_i_accept_w)
    ,.mem_i_valid_i(mem_i_valid_w)
    ,.mem_i_error_i(mem_i_error_w)
    ,.mem_i_inst_i(mem_i_inst_w)
    ,.intr_i(1'b0)
    ,.reset_vector_i(32'h80000000)
    ,.cpu_id_i('b0)
    ,.mem_d_addr_o(mem_d_addr_w)
    ,.mem_d_data_wr_o(mem_d_data_wr_w)
    ,.mem_d_rd_o(mem_d_rd_w)
    ,.mem_d_wr_o(mem_d_wr_w)
    ,.mem_d_cacheable_o(mem_d_cacheable_w)
    ,.mem_d_req_tag_o(mem_d_req_tag_w)
    ,.mem_d_invalidate_o(mem_d_invalidate_w)
    ,.mem_d_writeback_o(mem_d_writeback_w)
    ,.mem_d_flush_o(mem_d_flush_w)
    ,.mem_i_rd_o(mem_i_rd_w)
    ,.mem_i_flush_o(mem_i_flush_w)
    ,.mem_i_invalidate_o(mem_i_invalidate_w)
    ,.mem_i_pc_o(mem_i_pc_w)
);

tcm_mem u_mem
(
     .clk_i(clk)
    ,.rst_i(rst)
    ,.mem_i_rd_i(mem_i_rd_w)
    ,.mem_i_flush_i(mem_i_flush_w)
    ,.mem_i_invalidate_i(mem_i_invalidate_w)
    ,.mem_i_pc_i(mem_i_pc_w)
    ,.mem_d_addr_i(mem_d_addr_mem_w)
    ,.mem_d_data_wr_i(mem_d_data_wr_w)
    ,.mem_d_rd_i(mem_d_rd_w)
    ,.mem_d_wr_i(mem_d_wr_w)
    ,.mem_d_cacheable_i(mem_d_cacheable_w)
    ,.mem_d_req_tag_i(mem_d_req_tag_w)
    ,.mem_d_invalidate_i(mem_d_invalidate_w)
    ,.mem_d_writeback_i(mem_d_writeback_w)
    ,.mem_d_flush_i(mem_d_flush_w)
    ,.mem_i_accept_o(mem_i_accept_w)
    ,.mem_i_valid_o(mem_i_valid_w)
    ,.mem_i_error_o(mem_i_error_w)
    ,.mem_i_inst_o(mem_i_inst_w)
    ,.mem_d_data_rd_o(mem_d_data_rd_w)
    ,.mem_d_accept_o(mem_d_accept_w)
    ,.mem_d_ack_o(mem_d_ack_w)
    ,.mem_d_error_o(mem_d_error_w)
    ,.mem_d_resp_tag_o(mem_d_resp_tag_w)
);

endmodule
